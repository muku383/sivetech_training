package axi_test_pkg;
   
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   `include "axi_txn.sv";
   // `include "axi_cov.sv";
   `include "axi_drv.sv";
   `include "axi_mon.sv";
   `include "axi_seqr.sv";
   `include "axi_agent.sv";
   `include "axi_env.sv";
   `include "axi_seq.sv";
   `include "axi_test.sv";

endpackage
