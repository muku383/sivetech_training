
   //---------------------------------------------------------------------------
   // Typedef: ahb_sequencer
   //---------------------------------------------------------------------------

   typedef uvm_sequencer#(ahb_transaction) ahb_sequencer;
