`include "uvm_macros.svh"
   import uvm_pkg::*;
`timescale 1ps/1ps

`include "ahb_interfcae.sv"
`include "ahb_transaction.sv"
`include "ahb_reg_access_seq.sv"
`include "ahb_driver.sv"
`include "ahb_sequencer.sv"
`include "ahb_fc_subscriber.sv"
`include "ahb_monitor.sv"
`include "ahb_agent.sv"
`include "ahb_env.sv"
`include "ahb_base_test.sv"
`include "ahb_slave.sv"
`include "top.sv"
